module project_template(a,b,c);
       input a,b;
       output c;
       assign c=a|b;
endmodule
