module top(a,b,c);
    input a,b;
    output c;
    project_template project_template_inst(a,b,c);
endmodule