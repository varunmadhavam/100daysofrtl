module top(a,b,c);
    input a,b;
    output c;
    project_template dut(a,b,c);
endmodule